** sch_path: /foss/designs/Chipathon2024/ota-5t/xschem/ota-5t.sch
.subckt ota-5t Vp Vn Vout VDD VSS Ib
*.PININFO Vp:I Vn:I Vout:O VDD:B VSS:B Ib:I
XM2b Vout mirr VDD VDD sky130_fd_pr__pfet_01v8 L={l2} W={w2} nf={nf2} m=1
XM2a mirr mirr VDD VDD sky130_fd_pr__pfet_01v8 L={l2} W={w2} nf={nf2} m=1
XM1a mirr Vp tail VSS sky130_fd_pr__nfet_01v8_lvt L={l1} W={w1} nf={nf1} m=1
XM1b Vout Vn tail VSS sky130_fd_pr__nfet_01v8_lvt L={l1} W={w1} nf={nf1} m=1
XM0b tail Ib VSS VSS sky130_fd_pr__nfet_01v8_lvt L={l0} W={w0} nf={nf0} m=1
XM0a Ib Ib VSS VSS sky130_fd_pr__nfet_01v8_lvt L={l0} W={w0} nf={nf0} m=1
.ends
.end
