.param ib = 8.98e-05
.param cl = 1.68e-12
.param w0 = 371.57
.param l0 = 2.00
.param nf0 = 75.00
.param w1 = 185.79
.param l1 = 2.00
.param nf1 = 38.00
.param w2 = 2.76
.param l2 = 0.30
.param nf2 = 1.00
