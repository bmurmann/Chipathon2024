.param ib = 1.06e-05
.param cl = 1.78e-12
.param w0 = 23.23
.param l0 = 1.00
.param nf0 = 5.00
.param w1 = 5.83
.param l1 = 0.50
.param nf1 = 2.00
.param w2 = 1.13
.param l2 = 1.00
.param nf2 = 1.00
