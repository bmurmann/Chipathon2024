** sch_path: /foss/designs/Chipathon2024/techsweep_nfet_01v8_lvt.sch
**.subckt techsweep_nfet_01v8_lvt
vg g GND 0.9
vd d GND 0.9
vsb GND b {vbx}
XM1 d g GND b sky130_fd_pr__nfet_01v8_lvt L={lx} W={wx} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.param wx=5 lx=0.15 vbx=0
.dc vg 0 1.8 25m vd 0 1.8 25m
.control
option numdgt = 3
set wr_singlescale
set wr_vecnames

foreach l_val 0.15 0.16 0.17 0.18 0.19
+ 0.2 0.3 0.4 0.5 0.6 0.7 0.8 0.9 1 2 3
  alterparam lx = $l_val
  foreach vb_val 0 0.2 0.4
    alterparam vbx = $vb_val
    reset
    run
    wrdata techsweep_nfet_01v8_lvt.txt all
    destroy $curplot
    set appendwrite
  end
end
set appendwrite=0

alterparam lx = 0.15
alterparam vbx = 0
reset
op
showmod
show
write techsweep_nfet_01v8_lvt.raw
.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[capbd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[capbs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cdd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgb]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgd]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgg]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[cgs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[css]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gmbs]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[l]
.save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[vth]
.save b d g


**** end user architecture code
**.ends
.GLOBAL GND
.end
