** sch_path: /foss/designs/Chipathon2024/ota-5t/cace/templates/ota-5t_tb_noise.sch
**.subckt ota-5t_tb_noise
V0 VSS GND 0
V2 VDD GND {vdd}
E1 Vp net2 net1 GND 0.5
E2 Vn net2 net1 GND -0.5
Vdm net1 GND ac 1
Vcm net2 GND {vcm}
C2 Vout_buf GND {cl} m=1
x2 Vin_buf Vout_buf Vout_buf VDD VSS Ib ota-5t
Vibuf Vin_buf GND dc {vcm} ac 1
I1 VDD Ib {ib}
**** begin user architecture code


.lib {PDK_ROOT}/{PDK}/libs.tech/combined/sky130.lib.spice {corner}
.include {DUT_path}
.include /foss/designs/Chipathon2024/ota-5t/xschem/sizing_ota-5t.spice
.temp {temperature}




.control
    noise v(Vout_buf) Vibuf dec 20 1k 100e9
    setplot noise2
    let NOI = onoise_total/1e-6
    echo $&NOI > {simpath}/{filename}_{N}.data
    quit
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
