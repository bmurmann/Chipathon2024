.param ib = 3.67e-04
.param cl = 7.02e-12
.param w0 = 485.62
.param l0 = 0.60
.param nf0 = 98.00
.param w1 = 242.81
.param l1 = 0.60
.param nf1 = 49.00
.param w2 = 96.40
.param l2 = 0.60
.param nf2 = 20.00
