.param ib = 1e-05
.param cl = 1e-12
.param l0 = 1
.param l1 = 0.5
.param l2 = 1
.param w0 = 2.0
.param w1 = 20.0
.param w2 = 2.0
.param nf0 = 2
.param nf1 = 4
.param nf2 = 2
