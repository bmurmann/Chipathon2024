** sch_path: /foss/designs/Chipathon2024/techsweep_pfet_01v8.sch
**.subckt techsweep_pfet_01v8
Hn GND n vd 1
vg GND g DC 0.9 AC 1
vd GND d 0.9
vb GND b 0
XM1 d g GND b sky130_fd_pr__pfet_01v8 L={lx} W={wx} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.param wx=5 lx=0.15
.noise v(n) vg lin 1 1 1 1

.control
option numdgt = 3
set wr_singlescale
set wr_vecnames

compose l_vec  values 0.15 0.16 0.17 0.18 0.19
+ 0.2 0.3 0.4 0.5 0.6 0.7 0.8 0.9 1 2 3
compose vg_vec start= 0 stop=1.8  step=25m
compose vd_vec start= 0 stop=1.8  step=25m
compose vb_vec start= 0 stop=-0.4 step=-0.2

foreach var1 $&l_vec
  alterparam lx=$var1
  reset
  foreach var2 $&vg_vec
    alter vg $var2
    foreach var3 $&vd_vec
      alter vd $var3
      foreach var4 $&vb_vec
        alter vb $var4
        run
        wrdata techsweep_pfet_01v8.txt noise1.all
        destroy all
        set appendwrite
        unset set wr_vecnames
      end
    end
  end
end
unset appendwrite

alterparam lx=0.15
reset
op
show
write techsweep_pfet_01v8.raw
.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



.save @m.xm1.msky130_fd_pr__pfet_01v8[capbd]
.save @m.xm1.msky130_fd_pr__pfet_01v8[capbs]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cdd]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cgb]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cgd]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cgg]
.save @m.xm1.msky130_fd_pr__pfet_01v8[cgs]
.save @m.xm1.msky130_fd_pr__pfet_01v8[css]
.save @m.xm1.msky130_fd_pr__pfet_01v8[gds]
.save @m.xm1.msky130_fd_pr__pfet_01v8[gm]
.save @m.xm1.msky130_fd_pr__pfet_01v8[gmbs]
.save @m.xm1.msky130_fd_pr__pfet_01v8[id]
.save @m.xm1.msky130_fd_pr__pfet_01v8[l]
.save @m.xm1.msky130_fd_pr__pfet_01v8[vbs]
.save @m.xm1.msky130_fd_pr__pfet_01v8[vds]
.save @m.xm1.msky130_fd_pr__pfet_01v8[vgs]
.save @m.xm1.msky130_fd_pr__pfet_01v8[vth]
.save onoise.m.xm1.msky130_fd_pr__pfet_01v8.id
.save onoise.m.xm1.msky130_fd_pr__pfet_01v8.1overf
.save g d b n


**** end user architecture code
**.ends
.GLOBAL GND
.end
