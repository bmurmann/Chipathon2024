** sch_path: /foss/designs/chipathon/techsweep_nfet_01v8.sch
**.subckt techsweep_nfet_01v8
vg g GND 0.9
vd d GND 0.9
vb GND b {vbx}
XM1 d g GND b sky130_fd_pr__nfet_01v8 L={lx} W={wx} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.param wx=5 lx=0.15 vbx=0
.dc vg 0 1.8 25m vd 0 1.8 25m
.control
option numdgt = 3
set wr_singlescale
set wr_vecnames

foreach l_val 0.15 0.16 0.17 0.18 0.19
+ 0.2 0.3 0.4 0.5 0.6 0.7 0.8 0.9 1 2 3
  alterparam lx = $l_val
  foreach vb_val 0 0.2 0.4
    alterparam vbx = $vb_val
    reset
    run
   wrdata techsweep_nfet_01v8.txt all
    destroy $curplot
    set appendwrite
  end
end
set appendwrite=0

alterparam lx = 0.15
alterparam vbx = 0
reset
op
showmod
show
write techsweep_nfet_01v8.raw
.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



.save @m.xm1.msky130_fd_pr__nfet_01v8[capbd]
.save @m.xm1.msky130_fd_pr__nfet_01v8[capbs]
.save @m.xm1.msky130_fd_pr__nfet_01v8[cgg]
.save @m.xm1.msky130_fd_pr__nfet_01v8[gds]
.save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
.save @m.xm1.msky130_fd_pr__nfet_01v8[gmbs]
.save @m.xm1.msky130_fd_pr__nfet_01v8[id]
.save @m.xm1.msky130_fd_pr__nfet_01v8[l]
.save @m.xm1.msky130_fd_pr__nfet_01v8[vth]
.save b d g


**** end user architecture code
**.ends
.GLOBAL GND
.end
