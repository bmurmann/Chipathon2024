** sch_path: /foss/designs/chipathon/captest_nfet_01v8_lvt.sch
**.subckt captest_nfet_01v8_lvt
vg g GND dc 0.9 ac 1
vd d GND dc 0.9
vsb GND b {vsbx}
XM1 d g GND b sky130_fd_pr__nfet_01v8_lvt L={lx} W={wx} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.param wx=5 lx=0.15 vsbx=0
.param freq = 1Meg
.csparam freq = {freq}
.ac lin 1 {freq} {freq}

.control
run
print -im(vg#branch)/(2*PI*freq)
op
show
showmod m.XM1.msky130_fd_pr__nfet_01v8_lvt
.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
